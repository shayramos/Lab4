
module InterfaceAvalon (
	codecdata_bclk,
	codecdata_codecserialdata,
	codecdata_lrck);	

	output		codecdata_bclk;
	output		codecdata_codecserialdata;
	output		codecdata_lrck;
endmodule
