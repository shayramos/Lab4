
module InterfaceAvalon (
	codecdata_bclk,
	codecdata_codecserialdata,
	codecdata_lrck,
	clk_clk);	

	output		codecdata_bclk;
	output		codecdata_codecserialdata;
	output		codecdata_lrck;
	input		clk_clk;
endmodule
