
module InterfaceAvalon (
	clk_clk,
	codecdata_bclk,
	codecdata_codecserialdata,
	codecdata_lrck);	

	input		clk_clk;
	output		codecdata_bclk;
	output		codecdata_codecserialdata;
	output		codecdata_lrck;
endmodule
