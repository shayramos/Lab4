
module InterfaceAvalon (
	audioprocessor_0_conduit_end_bclk,
	audioprocessor_0_conduit_end_codecserialdata,
	audioprocessor_0_conduit_end_lrck,
	clk_clk);	

	output		audioprocessor_0_conduit_end_bclk;
	output		audioprocessor_0_conduit_end_codecserialdata;
	output		audioprocessor_0_conduit_end_lrck;
	input		clk_clk;
endmodule
